module Constant15(
	output [3:0] out
);

	assign out = 4'hF;
	
endmodule

module Constant4(
	output [31:0] out
);

	assign out = 32'h04;
	
endmodule

module Constant0(
	output out
);

	assign out = 1'b0;
	
endmodule